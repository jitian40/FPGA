module ip_core();

endmodule