module pll_simulation_test(
        input wire clk  //clock signal
);
endmodule  